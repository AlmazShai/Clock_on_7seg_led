`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:34:22 11/06/2020 
// Design Name: 
// Module Name:    Set_time 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Set_time(
    input key1,
    input key2,
    input key3,
    input key4,
    output [3:0] digit5,
    output [3:0] digit4,
    output [3:0] digit3,
    output [3:0] digit2,
    output [3:0] digit1,
    output [3:0] digit0,
    input clk,
    input reset
    );


endmodule
